* res_bcs corner
.lib "cornerRES.lib" mos_bcs
