* res_wcs corner
.lib "cornerRES.lib" mos_wcs
