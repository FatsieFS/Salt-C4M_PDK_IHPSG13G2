* lvmos_ff corner
.lib "cornerMOSlv.lib" mos_ff
