* hvmos_ff corner
.lib "cornerMOShv.lib" mos_ff
