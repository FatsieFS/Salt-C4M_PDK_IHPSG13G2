* hvmos_sf corner
.lib "cornerMOShv.lib" mos_sf
