* hvmos_tt corner
.lib "cornerMOShv.lib" mos_tt
