* res_typ corner
.lib "cornerRES.lib" mos_typ
