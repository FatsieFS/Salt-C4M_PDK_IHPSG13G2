* lvmos_sf corner
.lib "cornerMOSlv.lib" mos_sf
