* lvmos_fs corner
.lib "cornerMOSlv.lib" mos_fs
