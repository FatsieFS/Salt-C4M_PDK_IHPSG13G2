* hvmos_fs corner
.lib "cornerMOShv.lib" mos_fs
