* lvmos_tt corner
.lib "cornerMOSlv.lib" mos_tt
