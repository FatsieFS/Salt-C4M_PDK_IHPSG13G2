* lvmos_ss corner
.lib "cornerMOSlv.lib" mos_ss
