* hvmos_ss corner
.lib "cornerMOShv.lib" mos_ss
